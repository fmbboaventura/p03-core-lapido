module program_counter (
	input clk,    // Clock
	input [31:0] pc_in,

	output [31:0] pc_out
	
);

always @ (clk, pc_in, pc_out) begin 

end

endmodule